//testfile